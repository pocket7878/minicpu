`ifndef MINI_CPU_DEF_H
`define MINI_CPU_DEF_H

`define DATA_WIDTH 8
`define PROG_WIDTH 8

`endif