`include "def.svh"

module MINI_CPU_tb;
endmodule