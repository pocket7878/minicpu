`ifndef MINI_CPU_DEF_H
`define MINI_CPU_DEF_H

/**************************************
* [ 4bit op-code | 8bit immidiate ]
* <----------- Program ----------->
*                <--- register --->
***************************************/
`define DATA_WIDTH 8
`define OP_WIDTH 4
`define IM_WIDTH 8
`define PROG_WIDTH 12

`endif